module addi();

endmodule